package pack;
	
         import uvm_pkg::*;
	`include "uvm_macros.svh"

        `include "tb_config.sv"
        `include "xtn.sv"
        `include "seq.sv"
	`include "mon.sv"
	`include "drv.sv"
	`include "seqr.sv"
	`include "agt.sv"
	`include "sb.sv"
	`include "env.sv"
        `include "test.sv"

endpackage
        
        